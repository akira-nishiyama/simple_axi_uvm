package tb_simple_axi_uvm_test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import simple_axi_uvm_pkg::*;
    `include "tb_simple_axi_uvm_env.svh"
    `include "tb_simple_axi_uvm_sequence.svh"
    `include "tb_simple_axi_uvm_test.svh"

endpackage

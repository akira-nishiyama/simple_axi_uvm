package simple_axi_uvm_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "simple_axi_seq_item.svh"
    `include "simple_axi_master_sequencer.svh"
    `include "simple_axi_master_driver.svh"
    `include "simple_axi_master_monitor.svh"
    `include "simple_axi_master_agent.svh"
    `include "simple_axi_master_base_sequence.svh"
endpackage
